// pdp_11_const.vh
// Verilog include file with constants

`define DATA_MEMORY_SIZE 	16'hFFFF	//64K
`define FLASH_MEMORY_SIZE 	16'hFFFF	//64K